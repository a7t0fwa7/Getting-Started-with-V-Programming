//file: mod1/file3.v

module mod1

pub fn gday(){
	println('G\'Day Mother Fuckers from Mod1!!!!' )
}