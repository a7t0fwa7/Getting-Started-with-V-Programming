module mod1

pub const greet_msg = 'Greeting from mod1!'

/*
Accessing the constants of a module from another is a straightforward approach. 
You can access the constants of the module provided that they are marked as public using the pub keyword.

In our sample modulebasics project, let's consider the mod1 module with file1.v

In the preceding code, we have defined a constant named greet_msg in the mod1 module. Additionally, 
we marked the constant as public using the pub keyword.
*/
