module main

import mod1
import mod2

fn main() {
	mod1.hello()
	mod2.gday()
	println('Hello World!')
}
