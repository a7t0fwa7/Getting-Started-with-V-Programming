//file: mod2/file2.v

module mod2

pub fn gday(){
	println('Hello from mod2 mother fuckers!!')
}