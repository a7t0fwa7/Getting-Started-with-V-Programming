module main

fn main() {
	println('Hello World!')
}

/*Modular programming is the concept of logically grouping related functionalities together into modules and working with them. 
This approach enables you to wrap the related functionality into modules and allows you to import the required functionality that 
is available in those modules. 

V offers the concept of modular programming, allowing you to create and import modules that comprise code that is functionally or 
logically relevant in nature.
*/
