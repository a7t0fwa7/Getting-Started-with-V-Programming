module main

import mod1

fn main() {
	mod1.hello()
	//mod1.hello2()
}
